module Buffer(
	input in1,
	output out
);
	assign out = in1;
endmodule
