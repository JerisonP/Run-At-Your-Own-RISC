module NAND;
	logic 
